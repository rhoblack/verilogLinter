module test;
    `uvm_info("TEST", "Hello World", UVM_LOW)
endmodule
