`include "uvm_macros.svh"
import uvm_pkg::*;
module test;
    `uvm_info("TEST", "Hello World", UVM_LOW)
endmodule
